module ArithmeticLogicUnit(

);



endmodule


opcode 3 
000
001
010
011
100